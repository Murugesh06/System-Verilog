interface inf(input logic clk);
  logic rst;
  logic m;
  logic [3:0] count;
endinterface
