interface inf(input logic clk,rst,en);
  logic [3:0]addr;
  logic [7:0]data_in;
  logic [7:0]data_out;
endinterface
