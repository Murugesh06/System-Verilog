interface dff_if(input logic clk,rst);
  
  logic d;
  logic q;
  
endinterface
